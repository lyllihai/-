* test tran

VCC 1 0 3
R1 1 2 1000
C1 2 0 1e-5

.tran stop=0.04
.END